Bridge Rectifier

*declaring model
.MODEL DIO D( IS=1.8E-10 RS=2 BV=50.0 IBV=1e-4+ CJO=1e-12 M=0.333 N=2.06 TT=4.32e-9)

*resister between node 1 and 2
Rs 1 2 0.0011

*primary winding i.e. inductor
Lp 2 0 1mH
*secondary winding
Ls 3 4 1mH

*declaring diodes
D1 0 3 DIO
D2 3 5 DIO
D3 4 5 DIO
D4 0 4 DIO


*declaring coupling coefficients between inductors
Kps  Lp  Ls  1

*declaring capacitor
C1 5 0 0u

*load resister
RL 5 0 1K

*declaring sinusoidal voltage
v1 1 0 sin(0 16V 50)

*start the transient analysis
.tran 0.01m 40m

*control statement for simulation
.control

*run the simulation
run
*plot the curve between voltages on node 1 and 5
plot v(1) v(5)

*end of the control statement
.endc

*end of the netlist
.end
