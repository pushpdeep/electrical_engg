OPAMP BAND PASS FILTER

*iinclude the model file
.include UA741.txt

*declaring model
*  NON-INVERTING INPUT
*  | INVERTING INPUT
*  | | POSITIVE POWER SUPPLY
*  | | | NEGATIVE POWER SUPPLY
*  | | | | OUTPUT
*  | | | | |
X1 0 1 3 4 5 UA741

*declaring capacitor, try changing C1 = 0.47U
C1 2 6 2.2u
C2 1 5 0.01u
*declaring resisters try changing R2 = 6.8k
R1 1 2 1000K
R2 1 2 10K

Vcc 3 0 dc 15v
Vee 0 4 dc 15v

*declaring AC voltage source
V1 6 0 ac 4V

*start the AC analysis
.ac dec 10 2 200k
*.ac dec 10 0 50k

*control statement for simulation
.control
*run the simulation
run
*plot the output curve between voltage at node 5 and 6 in db i.e. output vs input
*plot db(v(5)/v(6))
*plot for output
plot db(v(5))
*end of the control statement
.endc
*end of the netlist
.end