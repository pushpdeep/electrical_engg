High pass filter with op amp 

*include the model file
.include UA741.txt

*declaring model
*  NON-INVERTING INPUT
*  | INVERTING INPUT
*  | | POSITIVE POWER SUPPLY
*  | | | NEGATIVE POWER SUPPLY
*  | | | | OUTPUT
*  | | | | |
X1 1 2 3 4 5 UA741
*declaring capacitor between nodes 1,0
C 1 6 0.1uF
*declaring resisters
R 1 0 1k
R1 2 0 1000k
R2 2 5 100k

Vcc 3 0 dc 15v
Vee 0 4 dc 15v

*declaring AC voltage source
V1 6 0 ac 4V

*start the AC analysis
.ac dec 10 150 1MEG
*control statement for simulation
.control
*run the simulation
run
*plot the output curve between voltage at node 5 and 6 in db
plot db(v(5))
*plot db(v(5)/v(6))
*end of the control statement
.endc
*end of the netlist
.end
