* Blue LED characterization

* SPICE model 
*Blue LED SPICE Model Data
.model BLUE D(IS = 2.659E-20 N = 2.63815 RS = 8.14349)
*Green LED SPICE Model Data
.model GREEN D(IS = 9.847E-17 N = 2.396 RS = 12.9816)
*Red LED SPICE Model Data
.model RED D (IS = 4.366E-25 N = 1.38167 RS = 3.00014)
*Yellow LED SPICE Model Data
.model YELLOW D (IS = 6.77E-22 N = 1.62 RS = 4.6779)
*White LED SPICE Model Data
.model WHITE D (IS = 1.2853E-15 N = 3.99 RS = 8.12296)

* Resistive Load
R1 1 2 100

* Diode
D1 2 0 BLUE

* Voltage Source
Vin 1 0 dc 5.0v

* DC analysis: Vin is swept from 0.0V to 6.0V in steps of 0.05V

.control 

dc Vin 0.0001 6 0.0001
run

plot -Vin#branch vs V(2) 
plot ln(-Vin#branch) vs V(2)

.endc

.end
