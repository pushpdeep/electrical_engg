Half Wave Rectifier


*declaring the model
.MODEL DIO D( IS=1.8E-10 RS=2 BV=50.0 IBV=1e-4+ CJO=1e-12 M=0.333 N=2.06 TT=4.32e-9)


*declaring the diode using the model 
D1 1 2 DIO
*declaring resister, try changing value of resister
RL 3 0 1K
*for adding capacitor, try changing value of capacitor
C1 3 0 0u
*declaring dc voltage source for measuring current
V2 2 3 dc 0V

*declaring sinusoidal voltage source
v1 1 0 sin(0 16V 50)

*start transient analysis
*.tran 0.0001ms 40ms
.tran 0.001ms 40ms

*start of control statement
.control
*run the simulation
run
*plotting input and output together
plot v(3), v(1)
*plot the current through diode
*plot i(V2)
*end of control statement
.endc

*end of netlist
.end

