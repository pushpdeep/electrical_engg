To Study Wave Shaping Circuit

*declaring model
.MODEL DIO D( IS=1.8E-10 RS=2 BV=50.0 IBV=1e-4+ CJO=1e-12 M=0.333 N=2.06 TT=4.32e-9)

*resister between nodes 1,2
Rs 1 2 1k

*declaring diode
D1 3 2 DIO

*declaring DC voltage source between nodes 3,0
V1 3 0 dc 3v

*declaring sinusoidal voltage 
Vs 1 0 sin(0 4V 1k)

*start the transient analysis
.tran 0.001m 2m

*control statement for simulation
.control
*run the simulation
run
*plot the output curve for voltage on node 1 and 2
plot v(1) V(2) 
*plot v(1) vs v(2)
*end of the control statement
.endc
*end of the netlist
.end
